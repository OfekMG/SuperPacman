// HartsMatrixBitMap File
// A two level bitmap. dosplaying harts on the screen Feb 2025
//(c) Technion IIT, Department of Electrical Engineering 2025

module HartsMatrixBitMap (
    input logic clk,
    input logic resetN,
    input logic [10:0] offsetX,// offset from top left  position
    input logic [10:0] offsetY,
    input logic InsideRectangle, //input that the pixel is within a bracket
    input logic random_hart,
    input logic collision_Smiley_Hart,
	 input logic collision_ghost_Hart,


    output logic drawingRequest, //output that the pixel should be dispalyed
    output logic [7:0] RGBout  //rgb value from the bitmap
 ) ;


localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32

localparam  int MAZE_NUMBER_OF__X_BITS = 5;  // 2^5 = 32, enough for 20 tiles
localparam  int MAZE_NUMBER_OF__Y_BITS = 4;  // 2^4 = 16, enough for 15 tiles

//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;
localparam  int MAZE_WIDTH_X = 1 << MAZE_NUMBER_OF__X_BITS ;
localparam  int MAZE_HEIGHT_Y = 1 << MAZE_NUMBER_OF__Y_BITS ;



logic [10:0] offsetX_LSB;
logic [10:0] offsetY_LSB;
logic [10:0] offsetX_MSB;
logic [10:0] offsetY_MSB;

// Get the pixel's coordinates WITHIN a 32x32 tile (lower 5 bits)
assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0]; 
assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0]; 

// Get the TILE's coordinates on the map grid (the higher bits)
assign offsetX_MSB  = offsetX[(TILE_NUMBER_OF_X_BITS + MAZE_NUMBER_OF__X_BITS - 1):TILE_NUMBER_OF_X_BITS];
assign offsetY_MSB  = offsetY[(TILE_NUMBER_OF_Y_BITS + MAZE_NUMBER_OF__Y_BITS - 1):TILE_NUMBER_OF_Y_BITS];



// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 8 *16
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares
// all numbers here are hard coded to simplify the understanding


logic [0:(MAZE_HEIGHT_Y-1)][0:(MAZE_WIDTH_X-1)] [3:0]  MazeBitMapMask ;
// The maze of the objects, a 16x32 array. Note: The visible portion is 15x20.
logic [0:15][0:31][3:0] MazeDefaultBitMapMask = '{
  // ROW 0: Top border
  '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
  // ROW 1
  '{1,0,0,0,1,0,0,0,0,1,0,0,0,0,1,0,0,1,1,0,0,0,0,1,0,0,0,0,0,0,0,1},
  // ROW 2
  '{1,0,1,0,1,0,1,1,0,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,0,1},
  // ROW 3
  '{1,0,1,0,0,0,0,1,0,0,0,1,0,0,0,1,0,1,1,0,0,1,0,0,0,1,0,0,0,1,0,1},
  // ROW 4
  '{1,0,1,1,1,0,1,1,0,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,0,1},
  // ROW 5
  '{1,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,1},
  // ROW 6
  '{1,1,0,1,1,0,1,1,1,0,1,1,1,0,1,1,1,1,1,1,1,0,1,1,1,0,1,1,0,1,1,1},
  // ROW 7
  '{1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1},
  // ROW 8
  '{1,1,1,0,1,1,0,1,1,1,1,0,1,1,0,1,1,1,1,0,1,1,0,1,1,1,1,0,1,1,1,1},
  // ROW 9
  '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1},
  // ROW 10
  '{1,0,1,1,1,0,1,1,0,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,1,0,1,0,1},
  // ROW 11
  '{1,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,1},
  // ROW 12
  '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,0,1,1,0,1,1,1},
  // ROW 13
  '{1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1},
  // ROW 14: Bottom border
  '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
  // ROW 15: Padding row
  '{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1}
};

 

 logic [3:0] [0:(TILE_HEIGHT_Y-1)][0:(TILE_WIDTH_X-1)] [7:0]  object_colors  = {{{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}},
{{{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}, // h3
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}}},
	{{{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}, // h2
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}}},
	{{{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}, // h1
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73},
	{8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73,8'h73}}}};
	
 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
    if(!resetN) begin
        RGBout <= 8'h00;
        MazeBitMapMask <= MazeDefaultBitMapMask; // copy default tabel
    end
    else begin
        RGBout <= TRANSPARENT_ENCODING; // default
        if (collision_Smiley_Hart && MazeBitMapMask[offsetY_MSB][offsetX_MSB] != 4'h1)
            MazeBitMapMask[offsetY_MSB][offsetX_MSB] <= 4'h00; // clear entry
        
        if (InsideRectangle == 1'b1)
            begin
                case (MazeBitMapMask[offsetY_MSB][offsetX_MSB])
                    4'h0: RGBout <= TRANSPARENT_ENCODING;
                    default: RGBout <= object_colors[MazeBitMapMask[offsetY_MSB][offsetX_MSB] - 1][offsetY_LSB][offsetX_LSB];
                endcase
            end
    end
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

