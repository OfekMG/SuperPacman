// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Feb 2025 
//(c) Technion IIT, Department of Electrical Engineering 2025 



module	HartsMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic random_hart,
					input logic collision_Smiley_Hart,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


localparam  int TILE_NUMBER_OF_X_BITS = 5;  // 2^5 = 32  everu object 
localparam  int TILE_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 

localparam  int MAZE_NUMBER_OF__X_BITS = 4;  // 2^4 = 16 / /the maze of the objects 
localparam  int MAZE_NUMBER_OF__Y_BITS = 3;  // 2^3 = 8 

//-----

localparam  int TILE_WIDTH_X = 1 << TILE_NUMBER_OF_X_BITS ;
localparam  int TILE_HEIGHT_Y = 1 <<  TILE_NUMBER_OF_Y_BITS ;
localparam  int MAZE_WIDTH_X = 1 << MAZE_NUMBER_OF__X_BITS ;
localparam  int MAZE_HEIGHT_Y = 1 << MAZE_NUMBER_OF__Y_BITS ;


 logic [10:0] offsetX_LSB  ;
 logic [10:0] offsetY_LSB  ; 
 logic [10:0] offsetX_MSB ;
 logic [10:0] offsetY_MSB  ;

 assign offsetX_LSB  = offsetX[(TILE_NUMBER_OF_X_BITS-1):0] ; // get lower bits 
 assign offsetY_LSB  = offsetY[(TILE_NUMBER_OF_Y_BITS-1):0] ; // get lower bits 
 assign offsetX_MSB  = offsetX[(TILE_NUMBER_OF_X_BITS + MAZE_NUMBER_OF__X_BITS -1 ):TILE_NUMBER_OF_X_BITS] ; // get higher bits 
 assign offsetY_MSB  = offsetY[(TILE_NUMBER_OF_Y_BITS + MAZE_NUMBER_OF__Y_BITS -1 ):TILE_NUMBER_OF_Y_BITS] ; // get higher bits 
 

 
// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 8 *16 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the understanding 


logic [0:(MAZE_HEIGHT_Y-1)][0:(MAZE_WIDTH_X-1)] [3:0]  MazeBitMapMask ;
// 2 - strongest
// 3 - mid
// 4 - broken almost
// 1 - normal  

logic [0:15][0:15][3:0] MazeDefaultBitMapMask = '{
    // Row 0
    {4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1},
    // Row 1
    {4'h1, 4'h2, 4'h2, 4'h1, 4'h2, 4'h2, 4'h2, 4'h2, 4'h2, 4'h2, 4'h2, 4'h1, 4'h2, 4'h2, 4'h2, 4'h1},
    // Row 2
    {4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h2, 4'h1},
    // Row 3
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h2, 4'h1},
    // Row 4
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h1, 4'h2, 4'h1},
    // Row 5
    {4'h1, 4'h2, 4'h2, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h2, 4'h1},
    // Row 6
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h2, 4'h1},
    // Row 7
    {4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1},
    // Row 8
    {4'h1, 4'h2, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h1, 4'h2, 4'h2, 4'h1},
    // Row 9
    {4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1},
    // Row 10
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h1, 4'h2, 4'h1},
    // Row 11
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h2, 4'h1},
    // Row 12
    {4'h1, 4'h2, 4'h2, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h2, 4'h1},
    // Row 13
    {4'h1, 4'h2, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h2, 4'h1},
    // Row 14
    {4'h1, 4'h2, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h2, 4'h1},
    // Row 15
    {4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1}
};

 

 logic [3:0] [0:(TILE_HEIGHT_Y-1)][0:(TILE_WIDTH_X-1)] [7:0]  object_colors  = {{
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h0e,8'h17,8'h9f,8'h9f,8'hff,8'hbf,8'h13,8'h12,8'h12,8'h12,8'h12,8'h13,8'hff,8'hdf,8'h13,8'h12,8'h12,8'h12,8'h12,8'h13,8'hff,8'hff,8'h9f,8'h9f,8'h12,8'h05,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h7f,8'hbf,8'h1f,8'h1b,8'h1b,8'h1f,8'hdf,8'h3f,8'h7f,8'h7f,8'h1f,8'h1b,8'h1b,8'h1f,8'hdf,8'h1f,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h17,8'h1b,8'h01,8'hff,8'h7b,8'h0d,8'h01,8'h7f,8'hff,8'h17,8'h01,8'h3f,8'h9f,8'h06,8'h06,8'hff,8'h1f,8'h05,8'h1b,8'hff,8'h1b,8'h01,8'h12,8'hbb,8'h32,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h7f,8'h1f,8'h13,8'h77,8'h0e,8'h01,8'h01,8'h01,8'h13,8'hdf,8'h3f,8'h13,8'h05,8'h01,8'h01,8'h06,8'h77,8'h7f,8'hbf,8'h0e,8'h01,8'h01,8'h01,8'h13,8'hff,8'h0e,8'h7f,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'hff,8'h1b,8'h13,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h06,8'h7f,8'h3f,8'h05,8'h01,8'h01,8'h05,8'h3f,8'h1f,8'h06,8'h01,8'h01,8'h01,8'h01,8'h01,8'h13,8'h0e,8'h7f,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'h9f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf4,8'h01,8'h17,8'h05,8'h01,8'h01,8'h01,8'h00,8'h05,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h0e,8'h01,8'h01,8'h01,8'hdf,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h13,8'hff,8'h17,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h00,8'h24,8'h13,8'h01,8'hfd,8'h20,8'h01,8'hff,8'h01,8'hf9,8'hfd,8'h24,8'h01,8'h01,8'h01,8'h01,8'h7f,8'hbf,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hff,8'h0e,8'h01,8'h01,8'h92,8'h01,8'h00,8'h01,8'h01,8'h0e,8'h64,8'h01,8'hf8,8'hf4,8'h01,8'h01,8'h24,8'hf8,8'hff,8'hf8,8'h00,8'h01,8'h12,8'hdf,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h13,8'hdf,8'h06,8'h01,8'h01,8'h05,8'h01,8'hf9,8'hff,8'h01,8'h01,8'h24,8'hf8,8'hf8,8'hf8,8'hf8,8'h01,8'h32,8'h01,8'h01,8'h01,8'h0e,8'hdf,8'h0e,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h05,8'h9f,8'h77,8'h01,8'h01,8'h05,8'hf9,8'hff,8'hfe,8'h6c,8'hf9,8'h00,8'hfc,8'hf8,8'hfc,8'hf8,8'hf4,8'h01,8'h01,8'hfc,8'h00,8'hbf,8'h3b,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h01,8'h13,8'h3f,8'h05,8'h01,8'hf8,8'hfe,8'hfe,8'hfc,8'h6c,8'h01,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'h24,8'hf8,8'h25,8'hdf,8'h13,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hdf,8'h32,8'h0e,8'h05,8'h13,8'hf8,8'hfd,8'hfd,8'hf8,8'hf8,8'h64,8'h00,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h01,8'hff,8'h6d,8'h0e,8'hdb,8'h1f,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h13,8'hdf,8'h7f,8'h0e,8'h01,8'hf9,8'h01,8'h01,8'h24,8'hf9,8'hf8,8'hf8,8'h01,8'h6d,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h05,8'h05,8'h00,8'h01,8'h01,8'h13,8'hdf,8'h9f,8'h06,8'h01,8'h01},
	{8'h01,8'h01,8'hdf,8'h9f,8'h06,8'h01,8'h01,8'h01,8'h01,8'h01,8'h64,8'h01,8'hf8,8'h24,8'h01,8'h24,8'hf8,8'hfc,8'h8c,8'h00,8'h01,8'hf8,8'h01,8'hfd,8'hf8,8'h01,8'h01,8'h0e,8'hff,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'hbf,8'hff,8'h0e,8'h01,8'h01,8'hd0,8'hfc,8'h24,8'hf9,8'h24,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h00,8'h20,8'h00,8'h01,8'h6c,8'hf8,8'hf8,8'h01,8'h01,8'h17,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h7f,8'hdf,8'h0e,8'h01,8'h20,8'hf8,8'h00,8'h00,8'hd5,8'hf8,8'hf8,8'h24,8'h64,8'h84,8'h00,8'hff,8'h24,8'hf4,8'hf8,8'h00,8'h64,8'h8c,8'h01,8'h12,8'hdf,8'h3f,8'h06,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'h9f,8'h32,8'h3f,8'h01,8'h71,8'h01,8'hf8,8'hf8,8'hf8,8'hf8,8'h24,8'h6c,8'hf8,8'hf8,8'hf8,8'h64,8'hff,8'h1f,8'h24,8'h01,8'h01,8'h1f,8'hbb,8'h37,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h01,8'h3f,8'h7f,8'h1f,8'h12,8'h6c,8'hf4,8'hf8,8'hf8,8'hf4,8'h05,8'hd0,8'hf8,8'hf8,8'hf8,8'hf4,8'hb0,8'hd4,8'h0e,8'h17,8'h3b,8'hdf,8'h13,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h0e,8'hdf,8'h0e,8'h65,8'h01,8'h01,8'h64,8'hf0,8'hf4,8'h64,8'h64,8'hf4,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h04,8'hf9,8'hf8,8'hd5,8'h9f,8'h9f,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hbf,8'h3b,8'h64,8'h01,8'h01,8'hf4,8'hf9,8'h2e,8'hf4,8'h01,8'h05,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'h00,8'h01,8'hf8,8'hf8,8'h01,8'h05,8'hdf,8'h13,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'h9f,8'h0e,8'h01,8'h01,8'h01,8'h24,8'hf8,8'h24,8'h01,8'hb5,8'h05,8'hf4,8'hf4,8'hf4,8'h8c,8'h01,8'h16,8'h01,8'h8c,8'h00,8'h05,8'h01,8'h13,8'hdf,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h3b,8'hdf,8'h13,8'h01,8'h01,8'h01,8'h01,8'h6d,8'h01,8'h01,8'hb6,8'hb5,8'h64,8'h01,8'h01,8'hf9,8'hfc,8'h00,8'h01,8'hfe,8'h01,8'h01,8'h01,8'h01,8'h01,8'h37,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'hff,8'h1f,8'h01,8'h01,8'h01,8'h01,8'h72,8'h71,8'h01,8'h01,8'h16,8'h05,8'h01,8'hf9,8'h01,8'hf5,8'hf8,8'h05,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h7f,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'h9f,8'h1f,8'h13,8'h13,8'h01,8'h01,8'h01,8'h01,8'h01,8'h12,8'hdf,8'h7f,8'h01,8'h64,8'h01,8'h01,8'hdf,8'hdf,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h13,8'h0e,8'h7f,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'h7f,8'h1b,8'h13,8'hff,8'h13,8'h05,8'h01,8'h05,8'h37,8'hdf,8'h3b,8'hdf,8'h12,8'h6d,8'h01,8'h12,8'hff,8'h3b,8'hdf,8'h37,8'h05,8'h01,8'h05,8'h13,8'hff,8'h0e,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h12,8'h1b,8'h01,8'h96,8'h32,8'h05,8'h05,8'h9f,8'hdf,8'h17,8'h01,8'h3b,8'hbf,8'h0e,8'h06,8'hff,8'h17,8'h01,8'h17,8'hff,8'h7f,8'h05,8'h0e,8'h76,8'h2e,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h05,8'h1b,8'h1b,8'h1b,8'h1f,8'h1f,8'h9f,8'h7f,8'h1f,8'h1b,8'h1b,8'h1f,8'hdf,8'hbf,8'h9f,8'h7f,8'h1f,8'h1b,8'h1b,8'h1f,8'hbf,8'h7f,8'h1f,8'h1b,8'h1b,8'h1b,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h0e,8'h12,8'h7a,8'h7f,8'hff,8'hbf,8'h12,8'h0e,8'h0e,8'h0e,8'h0e,8'h12,8'hdf,8'hbf,8'h12,8'h0e,8'h0e,8'h0e,8'h0e,8'h12,8'hff,8'hff,8'h7f,8'h7b,8'h0e,8'h05,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'hb6,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01}},
{{
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h01},
	{8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h05,8'h01},
	{8'h01,8'h01,8'h01,8'h37,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1b,8'h1b,8'h1b,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1b,8'h1b,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h0e,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h12,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'hff,8'hff,8'h1f,8'h1f,8'hff,8'hff,8'h1f,8'h1b,8'hff,8'h7f,8'h1f,8'h1f,8'hff,8'h7f,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h05,8'h17,8'h17,8'h12,8'h05,8'h01,8'h01,8'h01,8'h17,8'h17,8'h17,8'h05,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'hff,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h6d,8'h01,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'hda,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'hff,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'hff,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h05,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'hff,8'h05,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h01,8'h01,8'h01,8'hf4,8'hf4,8'hf4,8'hf4,8'h01,8'h01,8'h01,8'h01,8'hff,8'h01,8'h01,8'h01,8'h01,8'h13,8'h9f,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h17,8'h7f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hfd,8'hfe,8'hff,8'hfd,8'hf8,8'hf8,8'hf8,8'hf4,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hdf,8'h3f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h17,8'h1f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf9,8'hff,8'hff,8'hfd,8'hfc,8'hfc,8'hf8,8'hfc,8'hf8,8'hf4,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h1f,8'h05,8'h01,8'h00},
	{8'h01,8'h01,8'h37,8'h1f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'hfd,8'hff,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf4,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h1f,8'h05,8'h01,8'h00},
	{8'h01,8'h01,8'h17,8'hdf,8'h12,8'h01,8'h01,8'h00,8'h01,8'h01,8'hfc,8'hff,8'hfd,8'hf8,8'hf8,8'hf8,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'h01,8'h01,8'h01,8'h01,8'h01,8'h9f,8'h7f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'hff,8'h05,8'h01,8'h01,8'h00,8'h01,8'hf5,8'hfc,8'hf8,8'hf8,8'hf8,8'hf9,8'hd0,8'hf8,8'hd0,8'hfc,8'hf8,8'hf8,8'hf0,8'h24,8'h01,8'h00,8'h01,8'h01,8'h05,8'hff,8'h0e,8'h01,8'h00},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf5,8'hf4,8'h8c,8'h84,8'hf8,8'hf8,8'hf8,8'hf0,8'hf8,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hfc,8'hf8,8'h64,8'hf8,8'hf8,8'hf8,8'hf0,8'hf8,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'hff,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'h64,8'h8c,8'h8c,8'h60,8'hf8,8'hf8,8'hf8,8'hf0,8'h24,8'h01,8'h6d,8'h01,8'h01,8'h01,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h17,8'hff,8'h0e,8'h01,8'h00,8'h01,8'h01,8'h24,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf4,8'h00,8'h01,8'h01,8'h01,8'h01,8'h3f,8'h9f,8'h0d,8'h01,8'h01},
	{8'h01,8'h01,8'h12,8'h1f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf4,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h1f,8'h05,8'h00,8'h00},
	{8'h01,8'h01,8'h13,8'h1f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'h24,8'hf0,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h00,8'h01,8'h01,8'h01,8'h00,8'h01,8'hff,8'h1f,8'h05,8'h01,8'h00},
	{8'h01,8'h01,8'h16,8'h9f,8'h37,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h24,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'h04,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hbf,8'h7f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'hff,8'h0e,8'h01,8'h01,8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'h8c,8'hf4,8'hf4,8'hf4,8'hf4,8'hb0,8'h01,8'h01,8'h25,8'h01,8'h01,8'h01,8'h01,8'h01,8'h0e,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h25,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h01,8'h01,8'hff,8'h0e,8'h01,8'h00},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'hb6,8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h6d,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hda,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h1f,8'h3f,8'h01,8'h25,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h05,8'h01,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h1b,8'h1b,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h12,8'hbf,8'hdf,8'h7b,8'h05,8'h01,8'h01,8'h06,8'hbb,8'hdf,8'hdf,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h9f,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h7f,8'h9f,8'h7f,8'h7f,8'h7f,8'hff,8'hdf,8'h1f,8'h1f,8'hbf,8'hff,8'h9f,8'h7f,8'hff,8'h7f,8'h1f,8'h1f,8'hdf,8'hbf,8'h7f,8'h7f,8'h7f,8'h7f,8'h3f,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h12,8'h1b,8'h1b,8'h1f,8'h1f,8'h1b,8'h1b,8'h16,8'h32,8'h32,8'h16,8'h1b,8'h1b,8'h1b,8'h1b,8'h16,8'h32,8'h32,8'h16,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h16,8'h05,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h2d,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'hb6,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01}}},
	{{
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'hba,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h12,8'h13,8'h17,8'hff,8'hbf,8'h13,8'h12,8'h12,8'h12,8'h12,8'h13,8'h9f,8'h9f,8'h13,8'h12,8'h12,8'h12,8'h12,8'h13,8'hff,8'hff,8'h17,8'h13,8'h12,8'h01,8'h01,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h7f,8'h9f,8'h1f,8'h1b,8'h1b,8'h1f,8'hff,8'h7f,8'h7f,8'h7f,8'h1f,8'h1b,8'h1b,8'h1f,8'hff,8'h1f,8'h1b,8'h1b,8'h1b,8'h1b,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h01,8'hff,8'h77,8'h05,8'h01,8'h7f,8'hff,8'h17,8'h01,8'h7f,8'h9f,8'h06,8'h06,8'hff,8'h1f,8'h05,8'h1b,8'hff,8'h1b,8'h01,8'h12,8'hbb,8'h32,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h12,8'h1b,8'h13,8'h77,8'h0e,8'h01,8'h01,8'h01,8'h13,8'hff,8'h3f,8'h13,8'h06,8'h01,8'h01,8'h06,8'h13,8'h7f,8'hbf,8'h0e,8'h01,8'h01,8'h05,8'h13,8'hff,8'h0e,8'h3f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'hff,8'h1b,8'h13,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h06,8'h9f,8'hff,8'h05,8'h01,8'h00,8'h05,8'hdf,8'h7f,8'h06,8'h01,8'h01,8'h01,8'h01,8'h01,8'h13,8'h0e,8'h7f,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'h7f,8'h3b,8'h01,8'h01,8'h01,8'h01,8'hda,8'h01,8'h01,8'h01,8'h01,8'h05,8'h01,8'h01,8'h01,8'h2d,8'h05,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hdf,8'h12,8'h01,8'h01},
	{8'h01,8'hff,8'h0f,8'hff,8'h17,8'h01,8'h01,8'hdf,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h25,8'h01,8'h01,8'h7f,8'hbf,8'h06,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hff,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf4,8'hf4,8'hf4,8'hf4,8'h01,8'h01,8'h01,8'h01,8'hff,8'h01,8'h01,8'h01,8'h12,8'hbf,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h13,8'hbf,8'h06,8'h01,8'h01,8'h01,8'h01,8'h01,8'hf9,8'hfe,8'hff,8'hfd,8'hfc,8'hfc,8'hf8,8'hf4,8'h01,8'h01,8'h01,8'h01,8'h01,8'h12,8'hff,8'h0e,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h05,8'hbf,8'h36,8'h01,8'h01,8'h01,8'h01,8'hf9,8'hff,8'hff,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf4,8'h01,8'h01,8'h01,8'h01,8'hdf,8'h3b,8'h05,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h01,8'h13,8'hff,8'h05,8'h01,8'h01,8'hf9,8'hff,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf4,8'h01,8'h01,8'h05,8'hff,8'h13,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hdf,8'h32,8'h0e,8'h05,8'h01,8'h01,8'hfc,8'hff,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'h01,8'h01,8'h01,8'h0e,8'hdb,8'h77,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h13,8'hdf,8'h9f,8'h0e,8'h01,8'h01,8'h01,8'hf9,8'hfc,8'hfc,8'hfc,8'hfc,8'hf9,8'hd0,8'hf8,8'hac,8'hfc,8'hfc,8'hf8,8'hf0,8'h24,8'h01,8'h01,8'h01,8'h13,8'hdf,8'h9f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h7f,8'h9f,8'h06,8'h01,8'h01,8'h01,8'h01,8'hf8,8'hfc,8'hfc,8'hfc,8'hf4,8'hf5,8'hf4,8'h8c,8'h84,8'hf8,8'hfc,8'hf8,8'hf0,8'hf8,8'h01,8'h01,8'h01,8'h01,8'h0e,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h7f,8'hff,8'h0e,8'h01,8'h01,8'h01,8'h01,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hf8,8'h64,8'hfc,8'hfc,8'hf8,8'hf0,8'hf8,8'h01,8'h01,8'h01,8'h01,8'h17,8'hff,8'h12,8'h01,8'h01},
	{8'h01,8'h01,8'h0f,8'h9f,8'hdf,8'h0e,8'h01,8'h01,8'h01,8'hd4,8'hf8,8'hfc,8'hfc,8'hf8,8'h64,8'h8c,8'h8c,8'h64,8'hf8,8'hf8,8'hf8,8'hf0,8'h24,8'h01,8'h71,8'h01,8'h13,8'hdf,8'h3f,8'h06,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hbf,8'h33,8'hbf,8'h01,8'h01,8'h64,8'hf8,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf4,8'hf4,8'h00,8'h01,8'h01,8'h9f,8'hdf,8'h37,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h05,8'h3f,8'hdf,8'h05,8'h01,8'h01,8'hf4,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf8,8'h01,8'h01,8'h05,8'hff,8'h13,8'h05,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h0e,8'hdf,8'h0e,8'h01,8'h01,8'h01,8'h64,8'hf0,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h24,8'h01,8'h01,8'h01,8'hbf,8'h7b,8'h05,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1f,8'hbf,8'h1b,8'h01,8'h01,8'h01,8'h01,8'h01,8'h64,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'h24,8'h01,8'h01,8'h01,8'h01,8'h0e,8'hff,8'h12,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h9f,8'h9f,8'h05,8'h01,8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'hac,8'hf4,8'hf4,8'hf4,8'hf4,8'hb0,8'h01,8'h01,8'h6d,8'h05,8'h01,8'h01,8'h01,8'h13,8'hdf,8'h1f,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h3b,8'hdf,8'h12,8'h01,8'h01,8'h01,8'h25,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h37,8'hff,8'h0e,8'h01,8'h01},
	{8'h01,8'h01,8'hff,8'h1f,8'h01,8'h01,8'h01,8'h96,8'h01,8'hb6,8'h01,8'h01,8'h01,8'h01,8'h96,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h92,8'h01,8'h01,8'h01,8'h01,8'h7f,8'h32,8'h01,8'h01},
	{8'h01,8'h01,8'h76,8'h1f,8'h13,8'h13,8'h01,8'h01,8'h01,8'h01,8'h01,8'h12,8'hdf,8'h37,8'h01,8'hb6,8'h01,8'h01,8'hbf,8'hdf,8'h0e,8'h01,8'h01,8'h01,8'h01,8'h01,8'h13,8'h0e,8'h7f,8'h2e,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h13,8'hdf,8'h13,8'h05,8'h01,8'h05,8'h37,8'hdf,8'h3b,8'hbb,8'h96,8'h01,8'h01,8'h12,8'hbb,8'h3b,8'hdf,8'h36,8'h05,8'h01,8'h05,8'h13,8'hff,8'h0e,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h0e,8'h1b,8'h01,8'hbb,8'h32,8'h05,8'h05,8'h9f,8'hdf,8'h13,8'h01,8'h3f,8'hbf,8'h0e,8'h06,8'hff,8'h1b,8'h01,8'h17,8'hff,8'h7b,8'h05,8'h0e,8'h97,8'h0e,8'h01,8'h1b,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h1b,8'h1b,8'h1b,8'h1f,8'h1f,8'h9f,8'h9f,8'h1f,8'h1b,8'h1b,8'h1f,8'hdf,8'h9f,8'hbf,8'h7f,8'h1f,8'h1b,8'h1b,8'h1f,8'hbf,8'h3f,8'h1f,8'h1b,8'h1b,8'h1b,8'h32,8'h05,8'h01,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h0e,8'h0e,8'h13,8'hff,8'hbf,8'h0e,8'h0e,8'h0e,8'h0e,8'h0e,8'h12,8'h7f,8'h7f,8'h0e,8'h0e,8'h0e,8'h0e,8'h0e,8'h0e,8'hff,8'hff,8'h13,8'h0e,8'h0e,8'h01,8'h04,8'h01,8'h01},
	{8'h01,8'h01,8'h6d,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'hb6,8'h01},
	{8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01}}
	},
	{{
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h00,8'h00,8'h00,8'h05,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h01,8'hff,8'h00,8'h00,8'h01,8'h00,8'h00,8'hdb,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h00,8'h00,8'h00,8'h00,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf4,8'hf4,8'hf4,8'hf4,8'h00,8'h01,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h01,8'h00,8'h00,8'hf8,8'hfe,8'hff,8'hfe,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'hf8,8'hff,8'hff,8'hfd,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'hfd,8'hff,8'hfe,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hff,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf9,8'hd0,8'hf8,8'hd0,8'hfc,8'hf8,8'hf8,8'hf0,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'hf8,8'hfc,8'hf8,8'hf9,8'hf4,8'h8c,8'h64,8'hf8,8'hf8,8'hf8,8'hf0,8'hf8,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h01,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hfd,8'hf8,8'h64,8'hf8,8'hf8,8'hf8,8'hf0,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf4,8'hf8,8'hf8,8'hfc,8'hf8,8'h24,8'h8c,8'h8c,8'h20,8'hf8,8'hf8,8'hf8,8'hf0,8'h24,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf4,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf4,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hf0,8'hf4,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf4,8'hf0,8'hf4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h24,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'h00,8'h01,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hf4,8'hf4,8'hf4,8'hf4,8'hb0,8'h00,8'h00,8'h25,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h00,8'hb6,8'h00,8'h01,8'h00,8'h00,8'hb6,8'h01,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h2d,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h96,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}}}};
	
 
//
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		if (collision_Smiley_Hart)
			MazeBitMapMask[offsetY_MSB][offsetX_MSB] <= 4'h00;  // clear entry 
		
		if (InsideRectangle == 1'b1 )	
			begin 
		   	case (MazeBitMapMask[offsetY_MSB][offsetX_MSB])
					 4'h0 : RGBout <= TRANSPARENT_ENCODING ;
					 4'h1 : RGBout <= object_colors[random_hart][offsetY_LSB][offsetX_LSB]; 
					 4'h2 : RGBout <= object_colors[4'h1][offsetY_LSB][offsetX_LSB] ; 
					 4'h3 : RGBout <= object_colors[4'h2][offsetY_LSB][offsetX_LSB] ; 
					 4'h4 : RGBout <= object_colors[4'h3][offsetY_LSB][offsetX_LSB] ; 
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 

	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

